// 16 Bit AND Module with Structural Verilog by using the And1Bit module
module And16Bit(output[15:0] result,
					input[15:0] a, 
					input[15:0] b);

	And4Bit and1(result[3:0], a[3:0], b[3:0]);
	And4Bit and2(result[7:4], a[7:4], b[7:4]);
	And4Bit and3(result[11:8], a[11:8], b[11:8]);
	And4Bit and4(result[15:12], a[15:12], b[15:12]);

endmodule 