module CarryLookaheadLogic32Bit(output[1:0] c_ins, input[31:0] a, b, input c_in);
    // This is the logic for the SECOND LEVEL of the carry lookahead.

    // pi = ai XOR bi
    // gi = ai AND bi

    wire [31:0] p;
    wire [31:0] g;

    Xor32Bit x1(p, a, b);
    And32Bit a1(g, a, b);

    // c_ins[0] = g[15] + p[15] * g[14] + p[15] * p[14] * g[13] + ... + p[15] * ... * p[0] * c_in
    // c_ins[1] = g[31] + p[31] * g[30] + p[31] * p[30] * g[29] + ... + p[31] * ... * p[16] * c_ins[0]

    wire [15:0] p_g_0;

    and and1(p_g_0[0], p[15], g[14]);
    and and2(p_g_0[1], p[15], p[14], g[13]);
    and and3(p_g_0[2], p[15], p[14], p[13], g[12]);
    and and4(p_g_0[3], p[15], p[14], p[13], p[12], g[11]);
    and and5(p_g_0[4], p[15], p[14], p[13], p[12], p[11], g[10]);
    and and6(p_g_0[5], p[15], p[14], p[13], p[12], p[11], p[10], g[9]);
    and and7(p_g_0[6], p[15], p[14], p[13], p[12], p[11], p[10], p[9], g[8]);
    and and8(p_g_0[7], p[15], p[14], p[13], p[12], p[11], p[10], p[9], p[8], g[7]);
    and and9(p_g_0[8], p[15], p[14], p[13], p[12], p[11], p[10], p[9], p[8], p[7], g[6]);
    and and10(p_g_0[9], p[15], p[14], p[13], p[12], p[11], p[10], p[9], p[8], p[7], p[6], g[5]);
    and and11(p_g_0[10], p[15], p[14], p[13], p[12], p[11], p[10], p[9], p[8], p[7], p[6], p[5], g[4]);
    and and12(p_g_0[11], p[15], p[14], p[13], p[12], p[11], p[10], p[9], p[8], p[7], p[6], p[5], p[4], g[3]);
    and and13(p_g_0[12], p[15], p[14], p[13], p[12], p[11], p[10], p[9], p[8], p[7], p[6], p[5], p[4], p[3], g[2]);
    and and14(p_g_0[13], p[15], p[14], p[13], p[12], p[11], p[10], p[9], p[8], p[7], p[6], p[5], p[4], p[3], p[2], g[1]);
    and and15(p_g_0[14], p[15], p[14], p[13], p[12], p[11], p[10], p[9], p[8], p[7], p[6], p[5], p[4], p[3], p[2], p[1], g[0]);
    and and16(p_g_0[15], p[15], p[14], p[13], p[12], p[11], p[10], p[9], p[8], p[7], p[6], p[5], p[4], p[3], p[2], p[1], p[0], c_in);

    or or1(c_ins[0], g[15], p_g_0[0], p_g_0[1], p_g_0[2], p_g_0[3], p_g_0[4], p_g_0[5], p_g_0[6], p_g_0[7], p_g_0[8], p_g_0[9], p_g_0[10], p_g_0[11], p_g_0[12], p_g_0[13], p_g_0[14], p_g_0[15]);

    wire [15:0] p_g_1;

    and and17(p_g_1[0], p[31], g[30]);
    and and18(p_g_1[1], p[31], p[30], g[29]);
    and and19(p_g_1[2], p[31], p[30], p[29], g[28]);
    and and20(p_g_1[3], p[31], p[30], p[29], p[28], g[27]);
    and and21(p_g_1[4], p[31], p[30], p[29], p[28], p[27], g[26]);
    and and22(p_g_1[5], p[31], p[30], p[29], p[28], p[27], p[26], g[25]);
    and and23(p_g_1[6], p[31], p[30], p[29], p[28], p[27], p[26], p[25], g[24]);
    and and24(p_g_1[7], p[31], p[30], p[29], p[28], p[27], p[26], p[25], p[24], g[23]);
    and and25(p_g_1[8], p[31], p[30], p[29], p[28], p[27], p[26], p[25], p[24], p[23], g[22]);
    and and26(p_g_1[9], p[31], p[30], p[29], p[28], p[27], p[26], p[25], p[24], p[23], p[22], g[21]);
    and and27(p_g_1[10], p[31], p[30], p[29], p[28], p[27], p[26], p[25], p[24], p[23], p[22], p[21], g[20]);
    and and28(p_g_1[11], p[31], p[30], p[29], p[28], p[27], p[26], p[25], p[24], p[23], p[22], p[21], p[20], g[19]);
    and and29(p_g_1[12], p[31], p[30], p[29], p[28], p[27], p[26], p[25], p[24], p[23], p[22], p[21], p[20], p[19], g[18]);
    and and30(p_g_1[13], p[31], p[30], p[29], p[28], p[27], p[26], p[25], p[24], p[23], p[22], p[21], p[20], p[19], p[18], g[17]);
    and and31(p_g_1[14], p[31], p[30], p[29], p[28], p[27], p[26], p[25], p[24], p[23], p[22], p[21], p[20], p[19], p[18], p[17], g[16]);
    and and32(p_g_1[15], p[31], p[30], p[29], p[28], p[27], p[26], p[25], p[24], p[23], p[22], p[21], p[20], p[19], p[18], p[17], p[16], c_ins[0]);

    or or2(c_ins[1], g[31], p_g_1[0], p_g_1[1], p_g_1[2], p_g_1[3], p_g_1[4], p_g_1[5], p_g_1[6], p_g_1[7], p_g_1[8], p_g_1[9], p_g_1[10], p_g_1[11], p_g_1[12], p_g_1[13], p_g_1[14], p_g_1[15]);


endmodule 